module chorus #(
  parameter int width = 16
 ) (
  input logic clk,
  input logic rst,

  input logic signed [width-1:0] in_signal,
  output logic signed [width-1:0] out_signal

);
  

endmodule
