module softclip_lut #(
    parameter int width = 24
 ) (
    input logic signed [width-1:0] in_signal,
    output logic signed [width-1:0] out_signal
);

    logic [7:0] addr;
    assign addr = in_signal[width-1:width-8] + 8'd128;
    always_comb begin 
        case (addr)
            8'd  0 : out_signal = -24'sd8388607;
            8'd  1 : out_signal = -24'sd8386611;
            8'd  2 : out_signal = -24'sd8384521;
            8'd  3 : out_signal = -24'sd8382330;
            8'd  4 : out_signal = -24'sd8380035;
            8'd  5 : out_signal = -24'sd8377630;
            8'd  6 : out_signal = -24'sd8375111;
            8'd  7 : out_signal = -24'sd8372472;
            8'd  8 : out_signal = -24'sd8369707;
            8'd  9 : out_signal = -24'sd8366810;
            8'd 10 : out_signal = -24'sd8363775;
            8'd 11 : out_signal = -24'sd8360596;
            8'd 12 : out_signal = -24'sd8357265;
            8'd 13 : out_signal = -24'sd8353776;
            8'd 14 : out_signal = -24'sd8350121;
            8'd 15 : out_signal = -24'sd8346293;
            8'd 16 : out_signal = -24'sd8342282;
            8'd 17 : out_signal = -24'sd8338082;
            8'd 18 : out_signal = -24'sd8333682;
            8'd 19 : out_signal = -24'sd8329073;
            8'd 20 : out_signal = -24'sd8324245;
            8'd 21 : out_signal = -24'sd8319189;
            8'd 22 : out_signal = -24'sd8313894;
            8'd 23 : out_signal = -24'sd8308348;
            8'd 24 : out_signal = -24'sd8302540;
            8'd 25 : out_signal = -24'sd8296458;
            8'd 26 : out_signal = -24'sd8290088;
            8'd 27 : out_signal = -24'sd8283418;
            8'd 28 : out_signal = -24'sd8276433;
            8'd 29 : out_signal = -24'sd8269120;
            8'd 30 : out_signal = -24'sd8261462;
            8'd 31 : out_signal = -24'sd8253445;
            8'd 32 : out_signal = -24'sd8245051;
            8'd 33 : out_signal = -24'sd8236263;
            8'd 34 : out_signal = -24'sd8227063;
            8'd 35 : out_signal = -24'sd8217433;
            8'd 36 : out_signal = -24'sd8207352;
            8'd 37 : out_signal = -24'sd8196801;
            8'd 38 : out_signal = -24'sd8185758;
            8'd 39 : out_signal = -24'sd8174201;
            8'd 40 : out_signal = -24'sd8162106;
            8'd 41 : out_signal = -24'sd8149449;
            8'd 42 : out_signal = -24'sd8136206;
            8'd 43 : out_signal = -24'sd8122350;
            8'd 44 : out_signal = -24'sd8107854;
            8'd 45 : out_signal = -24'sd8092690;
            8'd 46 : out_signal = -24'sd8076827;
            8'd 47 : out_signal = -24'sd8060236;
            8'd 48 : out_signal = -24'sd8042885;
            8'd 49 : out_signal = -24'sd8024740;
            8'd 50 : out_signal = -24'sd8005767;
            8'd 51 : out_signal = -24'sd7985930;
            8'd 52 : out_signal = -24'sd7965193;
            8'd 53 : out_signal = -24'sd7943516;
            8'd 54 : out_signal = -24'sd7920861;
            8'd 55 : out_signal = -24'sd7897186;
            8'd 56 : out_signal = -24'sd7872448;
            8'd 57 : out_signal = -24'sd7846603;
            8'd 58 : out_signal = -24'sd7819605;
            8'd 59 : out_signal = -24'sd7791408;
            8'd 60 : out_signal = -24'sd7761963;
            8'd 61 : out_signal = -24'sd7731218;
            8'd 62 : out_signal = -24'sd7699124;
            8'd 63 : out_signal = -24'sd7665625;
            8'd 64 : out_signal = -24'sd7630669;
            8'd 65 : out_signal = -24'sd7594197;
            8'd 66 : out_signal = -24'sd7556152;
            8'd 67 : out_signal = -24'sd7516474;
            8'd 68 : out_signal = -24'sd7475103;
            8'd 69 : out_signal = -24'sd7431977;
            8'd 70 : out_signal = -24'sd7387031;
            8'd 71 : out_signal = -24'sd7340201;
            8'd 72 : out_signal = -24'sd7291420;
            8'd 73 : out_signal = -24'sd7240620;
            8'd 74 : out_signal = -24'sd7187734;
            8'd 75 : out_signal = -24'sd7132692;
            8'd 76 : out_signal = -24'sd7075422;
            8'd 77 : out_signal = -24'sd7015855;
            8'd 78 : out_signal = -24'sd6953919;
            8'd 79 : out_signal = -24'sd6889540;
            8'd 80 : out_signal = -24'sd6822648;
            8'd 81 : out_signal = -24'sd6753170;
            8'd 82 : out_signal = -24'sd6681033;
            8'd 83 : out_signal = -24'sd6606167;
            8'd 84 : out_signal = -24'sd6528499;
            8'd 85 : out_signal = -24'sd6447961;
            8'd 86 : out_signal = -24'sd6364483;
            8'd 87 : out_signal = -24'sd6277998;
            8'd 88 : out_signal = -24'sd6188441;
            8'd 89 : out_signal = -24'sd6095749;
            8'd 90 : out_signal = -24'sd5999862;
            8'd 91 : out_signal = -24'sd5900722;
            8'd 92 : out_signal = -24'sd5798276;
            8'd 93 : out_signal = -24'sd5692473;
            8'd 94 : out_signal = -24'sd5583268;
            8'd 95 : out_signal = -24'sd5470621;
            8'd 96 : out_signal = -24'sd5354494;
            8'd 97 : out_signal = -24'sd5234859;
            8'd 98 : out_signal = -24'sd5111690;
            8'd 99 : out_signal = -24'sd4984971;
            8'd100 : out_signal = -24'sd4854691;
            8'd101 : out_signal = -24'sd4720847;
            8'd102 : out_signal = -24'sd4583443;
            8'd103 : out_signal = -24'sd4442493;
            8'd104 : out_signal = -24'sd4298018;
            8'd105 : out_signal = -24'sd4150050;
            8'd106 : out_signal = -24'sd3998627;
            8'd107 : out_signal = -24'sd3843801;
            8'd108 : out_signal = -24'sd3685631;
            8'd109 : out_signal = -24'sd3524187;
            8'd110 : out_signal = -24'sd3359548;
            8'd111 : out_signal = -24'sd3191805;
            8'd112 : out_signal = -24'sd3021059;
            8'd113 : out_signal = -24'sd2847421;
            8'd114 : out_signal = -24'sd2671013;
            8'd115 : out_signal = -24'sd2491966;
            8'd116 : out_signal = -24'sd2310421;
            8'd117 : out_signal = -24'sd2126529;
            8'd118 : out_signal = -24'sd1940450;
            8'd119 : out_signal = -24'sd1752352;
            8'd120 : out_signal = -24'sd1562414;
            8'd121 : out_signal = -24'sd1370818;
            8'd122 : out_signal = -24'sd1177757;
            8'd123 : out_signal = -24'sd983428;
            8'd124 : out_signal = -24'sd788033;
            8'd125 : out_signal = -24'sd591780;
            8'd126 : out_signal = -24'sd394881;
            8'd127 : out_signal = -24'sd197549;
            8'd128 : out_signal = 24'sd0;
            8'd129 : out_signal = 24'sd197549;
            8'd130 : out_signal = 24'sd394881;
            8'd131 : out_signal = 24'sd591780;
            8'd132 : out_signal = 24'sd788033;
            8'd133 : out_signal = 24'sd983428;
            8'd134 : out_signal = 24'sd1177757;
            8'd135 : out_signal = 24'sd1370818;
            8'd136 : out_signal = 24'sd1562414;
            8'd137 : out_signal = 24'sd1752352;
            8'd138 : out_signal = 24'sd1940450;
            8'd139 : out_signal = 24'sd2126529;
            8'd140 : out_signal = 24'sd2310421;
            8'd141 : out_signal = 24'sd2491966;
            8'd142 : out_signal = 24'sd2671013;
            8'd143 : out_signal = 24'sd2847421;
            8'd144 : out_signal = 24'sd3021059;
            8'd145 : out_signal = 24'sd3191805;
            8'd146 : out_signal = 24'sd3359548;
            8'd147 : out_signal = 24'sd3524187;
            8'd148 : out_signal = 24'sd3685631;
            8'd149 : out_signal = 24'sd3843801;
            8'd150 : out_signal = 24'sd3998627;
            8'd151 : out_signal = 24'sd4150050;
            8'd152 : out_signal = 24'sd4298018;
            8'd153 : out_signal = 24'sd4442493;
            8'd154 : out_signal = 24'sd4583443;
            8'd155 : out_signal = 24'sd4720847;
            8'd156 : out_signal = 24'sd4854691;
            8'd157 : out_signal = 24'sd4984971;
            8'd158 : out_signal = 24'sd5111690;
            8'd159 : out_signal = 24'sd5234859;
            8'd160 : out_signal = 24'sd5354494;
            8'd161 : out_signal = 24'sd5470621;
            8'd162 : out_signal = 24'sd5583268;
            8'd163 : out_signal = 24'sd5692473;
            8'd164 : out_signal = 24'sd5798276;
            8'd165 : out_signal = 24'sd5900722;
            8'd166 : out_signal = 24'sd5999862;
            8'd167 : out_signal = 24'sd6095749;
            8'd168 : out_signal = 24'sd6188441;
            8'd169 : out_signal = 24'sd6277998;
            8'd170 : out_signal = 24'sd6364483;
            8'd171 : out_signal = 24'sd6447961;
            8'd172 : out_signal = 24'sd6528499;
            8'd173 : out_signal = 24'sd6606167;
            8'd174 : out_signal = 24'sd6681033;
            8'd175 : out_signal = 24'sd6753170;
            8'd176 : out_signal = 24'sd6822648;
            8'd177 : out_signal = 24'sd6889540;
            8'd178 : out_signal = 24'sd6953919;
            8'd179 : out_signal = 24'sd7015855;
            8'd180 : out_signal = 24'sd7075422;
            8'd181 : out_signal = 24'sd7132692;
            8'd182 : out_signal = 24'sd7187734;
            8'd183 : out_signal = 24'sd7240620;
            8'd184 : out_signal = 24'sd7291420;
            8'd185 : out_signal = 24'sd7340201;
            8'd186 : out_signal = 24'sd7387031;
            8'd187 : out_signal = 24'sd7431977;
            8'd188 : out_signal = 24'sd7475103;
            8'd189 : out_signal = 24'sd7516474;
            8'd190 : out_signal = 24'sd7556152;
            8'd191 : out_signal = 24'sd7594197;
            8'd192 : out_signal = 24'sd7630669;
            8'd193 : out_signal = 24'sd7665625;
            8'd194 : out_signal = 24'sd7699124;
            8'd195 : out_signal = 24'sd7731218;
            8'd196 : out_signal = 24'sd7761963;
            8'd197 : out_signal = 24'sd7791408;
            8'd198 : out_signal = 24'sd7819605;
            8'd199 : out_signal = 24'sd7846603;
            8'd200 : out_signal = 24'sd7872448;
            8'd201 : out_signal = 24'sd7897186;
            8'd202 : out_signal = 24'sd7920861;
            8'd203 : out_signal = 24'sd7943516;
            8'd204 : out_signal = 24'sd7965193;
            8'd205 : out_signal = 24'sd7985930;
            8'd206 : out_signal = 24'sd8005767;
            8'd207 : out_signal = 24'sd8024740;
            8'd208 : out_signal = 24'sd8042885;
            8'd209 : out_signal = 24'sd8060236;
            8'd210 : out_signal = 24'sd8076827;
            8'd211 : out_signal = 24'sd8092690;
            8'd212 : out_signal = 24'sd8107854;
            8'd213 : out_signal = 24'sd8122350;
            8'd214 : out_signal = 24'sd8136206;
            8'd215 : out_signal = 24'sd8149449;
            8'd216 : out_signal = 24'sd8162106;
            8'd217 : out_signal = 24'sd8174201;
            8'd218 : out_signal = 24'sd8185758;
            8'd219 : out_signal = 24'sd8196801;
            8'd220 : out_signal = 24'sd8207352;
            8'd221 : out_signal = 24'sd8217433;
            8'd222 : out_signal = 24'sd8227063;
            8'd223 : out_signal = 24'sd8236263;
            8'd224 : out_signal = 24'sd8245051;
            8'd225 : out_signal = 24'sd8253445;
            8'd226 : out_signal = 24'sd8261462;
            8'd227 : out_signal = 24'sd8269120;
            8'd228 : out_signal = 24'sd8276433;
            8'd229 : out_signal = 24'sd8283418;
            8'd230 : out_signal = 24'sd8290088;
            8'd231 : out_signal = 24'sd8296458;
            8'd232 : out_signal = 24'sd8302540;
            8'd233 : out_signal = 24'sd8308348;
            8'd234 : out_signal = 24'sd8313894;
            8'd235 : out_signal = 24'sd8319189;
            8'd236 : out_signal = 24'sd8324245;
            8'd237 : out_signal = 24'sd8329073;
            8'd238 : out_signal = 24'sd8333682;
            8'd239 : out_signal = 24'sd8338082;
            8'd240 : out_signal = 24'sd8342282;
            8'd241 : out_signal = 24'sd8346293;
            8'd242 : out_signal = 24'sd8350121;
            8'd243 : out_signal = 24'sd8353776;
            8'd244 : out_signal = 24'sd8357265;
            8'd245 : out_signal = 24'sd8360596;
            8'd246 : out_signal = 24'sd8363775;
            8'd247 : out_signal = 24'sd8366810;
            8'd248 : out_signal = 24'sd8369707;
            8'd249 : out_signal = 24'sd8372472;
            8'd250 : out_signal = 24'sd8375111;
            8'd251 : out_signal = 24'sd8377630;
            8'd252 : out_signal = 24'sd8380035;
            8'd253 : out_signal = 24'sd8382330;
            8'd254 : out_signal = 24'sd8384521;
            8'd255 : out_signal = 24'sd8386611;
            default: out_signal = in_signal;
        endcase
    end

endmodule
            
