module softclip_lut (
    input logic signed [15:0] in_signal,
    output logic signed [15:0] out_signal
);


    logic [7:0] addr;
    assign addr = in_signal[15:8] + 8'd128;
    always_comb begin 
        case (addr)
            8'd  0 : out_signal = -16'sd32767;
            8'd  1 : out_signal = -16'sd32759;
            8'd  2 : out_signal = -16'sd32751;
            8'd  3 : out_signal = -16'sd32742;
            8'd  4 : out_signal = -16'sd32734;
            8'd  5 : out_signal = -16'sd32724;
            8'd  6 : out_signal = -16'sd32714;
            8'd  7 : out_signal = -16'sd32704;
            8'd  8 : out_signal = -16'sd32693;
            8'd  9 : out_signal = -16'sd32682;
            8'd 10 : out_signal = -16'sd32670;
            8'd 11 : out_signal = -16'sd32658;
            8'd 12 : out_signal = -16'sd32645;
            8'd 13 : out_signal = -16'sd32631;
            8'd 14 : out_signal = -16'sd32617;
            8'd 15 : out_signal = -16'sd32602;
            8'd 16 : out_signal = -16'sd32586;
            8'd 17 : out_signal = -16'sd32570;
            8'd 18 : out_signal = -16'sd32552;
            8'd 19 : out_signal = -16'sd32534;
            8'd 20 : out_signal = -16'sd32516;
            8'd 21 : out_signal = -16'sd32496;
            8'd 22 : out_signal = -16'sd32475;
            8'd 23 : out_signal = -16'sd32453;
            8'd 24 : out_signal = -16'sd32431;
            8'd 25 : out_signal = -16'sd32407;
            8'd 26 : out_signal = -16'sd32382;
            8'd 27 : out_signal = -16'sd32356;
            8'd 28 : out_signal = -16'sd32329;
            8'd 29 : out_signal = -16'sd32300;
            8'd 30 : out_signal = -16'sd32270;
            8'd 31 : out_signal = -16'sd32239;
            8'd 32 : out_signal = -16'sd32206;
            8'd 33 : out_signal = -16'sd32172;
            8'd 34 : out_signal = -16'sd32136;
            8'd 35 : out_signal = -16'sd32098;
            8'd 36 : out_signal = -16'sd32059;
            8'd 37 : out_signal = -16'sd32018;
            8'd 38 : out_signal = -16'sd31975;
            8'd 39 : out_signal = -16'sd31930;
            8'd 40 : out_signal = -16'sd31882;
            8'd 41 : out_signal = -16'sd31833;
            8'd 42 : out_signal = -16'sd31781;
            8'd 43 : out_signal = -16'sd31727;
            8'd 44 : out_signal = -16'sd31670;
            8'd 45 : out_signal = -16'sd31611;
            8'd 46 : out_signal = -16'sd31549;
            8'd 47 : out_signal = -16'sd31484;
            8'd 48 : out_signal = -16'sd31417;
            8'd 49 : out_signal = -16'sd31346;
            8'd 50 : out_signal = -16'sd31272;
            8'd 51 : out_signal = -16'sd31194;
            8'd 52 : out_signal = -16'sd31113;
            8'd 53 : out_signal = -16'sd31028;
            8'd 54 : out_signal = -16'sd30940;
            8'd 55 : out_signal = -16'sd30847;
            8'd 56 : out_signal = -16'sd30751;
            8'd 57 : out_signal = -16'sd30650;
            8'd 58 : out_signal = -16'sd30544;
            8'd 59 : out_signal = -16'sd30434;
            8'd 60 : out_signal = -16'sd30319;
            8'd 61 : out_signal = -16'sd30199;
            8'd 62 : out_signal = -16'sd30074;
            8'd 63 : out_signal = -16'sd29943;
            8'd 64 : out_signal = -16'sd29806;
            8'd 65 : out_signal = -16'sd29664;
            8'd 66 : out_signal = -16'sd29515;
            8'd 67 : out_signal = -16'sd29360;
            8'd 68 : out_signal = -16'sd29199;
            8'd 69 : out_signal = -16'sd29030;
            8'd 70 : out_signal = -16'sd28855;
            8'd 71 : out_signal = -16'sd28672;
            8'd 72 : out_signal = -16'sd28481;
            8'd 73 : out_signal = -16'sd28283;
            8'd 74 : out_signal = -16'sd28076;
            8'd 75 : out_signal = -16'sd27861;
            8'd 76 : out_signal = -16'sd27638;
            8'd 77 : out_signal = -16'sd27405;
            8'd 78 : out_signal = -16'sd27163;
            8'd 79 : out_signal = -16'sd26911;
            8'd 80 : out_signal = -16'sd26650;
            8'd 81 : out_signal = -16'sd26379;
            8'd 82 : out_signal = -16'sd26097;
            8'd 83 : out_signal = -16'sd25805;
            8'd 84 : out_signal = -16'sd25501;
            8'd 85 : out_signal = -16'sd25187;
            8'd 86 : out_signal = -16'sd24861;
            8'd 87 : out_signal = -16'sd24523;
            8'd 88 : out_signal = -16'sd24173;
            8'd 89 : out_signal = -16'sd23811;
            8'd 90 : out_signal = -16'sd23436;
            8'd 91 : out_signal = -16'sd23049;
            8'd 92 : out_signal = -16'sd22649;
            8'd 93 : out_signal = -16'sd22236;
            8'd 94 : out_signal = -16'sd21809;
            8'd 95 : out_signal = -16'sd21369;
            8'd 96 : out_signal = -16'sd20915;
            8'd 97 : out_signal = -16'sd20448;
            8'd 98 : out_signal = -16'sd19967;
            8'd 99 : out_signal = -16'sd19472;
            8'd100 : out_signal = -16'sd18963;
            8'd101 : out_signal = -16'sd18440;
            8'd102 : out_signal = -16'sd17904;
            8'd103 : out_signal = -16'sd17353;
            8'd104 : out_signal = -16'sd16789;
            8'd105 : out_signal = -16'sd16211;
            8'd106 : out_signal = -16'sd15619;
            8'd107 : out_signal = -16'sd15014;
            8'd108 : out_signal = -16'sd14397;
            8'd109 : out_signal = -16'sd13766;
            8'd110 : out_signal = -16'sd13123;
            8'd111 : out_signal = -16'sd12468;
            8'd112 : out_signal = -16'sd11801;
            8'd113 : out_signal = -16'sd11122;
            8'd114 : out_signal = -16'sd10433;
            8'd115 : out_signal = -16'sd9734;
            8'd116 : out_signal = -16'sd9025;
            8'd117 : out_signal = -16'sd8306;
            8'd118 : out_signal = -16'sd7580;
            8'd119 : out_signal = -16'sd6845;
            8'd120 : out_signal = -16'sd6103;
            8'd121 : out_signal = -16'sd5355;
            8'd122 : out_signal = -16'sd4600;
            8'd123 : out_signal = -16'sd3841;
            8'd124 : out_signal = -16'sd3078;
            8'd125 : out_signal = -16'sd2312;
            8'd126 : out_signal = -16'sd1542;
            8'd127 : out_signal = -16'sd772;
            8'd128 : out_signal = 16'sd0;
            8'd129 : out_signal = 16'sd772;
            8'd130 : out_signal = 16'sd1542;
            8'd131 : out_signal = 16'sd2312;
            8'd132 : out_signal = 16'sd3078;
            8'd133 : out_signal = 16'sd3841;
            8'd134 : out_signal = 16'sd4600;
            8'd135 : out_signal = 16'sd5355;
            8'd136 : out_signal = 16'sd6103;
            8'd137 : out_signal = 16'sd6845;
            8'd138 : out_signal = 16'sd7580;
            8'd139 : out_signal = 16'sd8306;
            8'd140 : out_signal = 16'sd9025;
            8'd141 : out_signal = 16'sd9734;
            8'd142 : out_signal = 16'sd10433;
            8'd143 : out_signal = 16'sd11122;
            8'd144 : out_signal = 16'sd11801;
            8'd145 : out_signal = 16'sd12468;
            8'd146 : out_signal = 16'sd13123;
            8'd147 : out_signal = 16'sd13766;
            8'd148 : out_signal = 16'sd14397;
            8'd149 : out_signal = 16'sd15014;
            8'd150 : out_signal = 16'sd15619;
            8'd151 : out_signal = 16'sd16211;
            8'd152 : out_signal = 16'sd16789;
            8'd153 : out_signal = 16'sd17353;
            8'd154 : out_signal = 16'sd17904;
            8'd155 : out_signal = 16'sd18440;
            8'd156 : out_signal = 16'sd18963;
            8'd157 : out_signal = 16'sd19472;
            8'd158 : out_signal = 16'sd19967;
            8'd159 : out_signal = 16'sd20448;
            8'd160 : out_signal = 16'sd20915;
            8'd161 : out_signal = 16'sd21369;
            8'd162 : out_signal = 16'sd21809;
            8'd163 : out_signal = 16'sd22236;
            8'd164 : out_signal = 16'sd22649;
            8'd165 : out_signal = 16'sd23049;
            8'd166 : out_signal = 16'sd23436;
            8'd167 : out_signal = 16'sd23811;
            8'd168 : out_signal = 16'sd24173;
            8'd169 : out_signal = 16'sd24523;
            8'd170 : out_signal = 16'sd24861;
            8'd171 : out_signal = 16'sd25187;
            8'd172 : out_signal = 16'sd25501;
            8'd173 : out_signal = 16'sd25805;
            8'd174 : out_signal = 16'sd26097;
            8'd175 : out_signal = 16'sd26379;
            8'd176 : out_signal = 16'sd26650;
            8'd177 : out_signal = 16'sd26911;
            8'd178 : out_signal = 16'sd27163;
            8'd179 : out_signal = 16'sd27405;
            8'd180 : out_signal = 16'sd27638;
            8'd181 : out_signal = 16'sd27861;
            8'd182 : out_signal = 16'sd28076;
            8'd183 : out_signal = 16'sd28283;
            8'd184 : out_signal = 16'sd28481;
            8'd185 : out_signal = 16'sd28672;
            8'd186 : out_signal = 16'sd28855;
            8'd187 : out_signal = 16'sd29030;
            8'd188 : out_signal = 16'sd29199;
            8'd189 : out_signal = 16'sd29360;
            8'd190 : out_signal = 16'sd29515;
            8'd191 : out_signal = 16'sd29664;
            8'd192 : out_signal = 16'sd29806;
            8'd193 : out_signal = 16'sd29943;
            8'd194 : out_signal = 16'sd30074;
            8'd195 : out_signal = 16'sd30199;
            8'd196 : out_signal = 16'sd30319;
            8'd197 : out_signal = 16'sd30434;
            8'd198 : out_signal = 16'sd30544;
            8'd199 : out_signal = 16'sd30650;
            8'd200 : out_signal = 16'sd30751;
            8'd201 : out_signal = 16'sd30847;
            8'd202 : out_signal = 16'sd30940;
            8'd203 : out_signal = 16'sd31028;
            8'd204 : out_signal = 16'sd31113;
            8'd205 : out_signal = 16'sd31194;
            8'd206 : out_signal = 16'sd31272;
            8'd207 : out_signal = 16'sd31346;
            8'd208 : out_signal = 16'sd31417;
            8'd209 : out_signal = 16'sd31484;
            8'd210 : out_signal = 16'sd31549;
            8'd211 : out_signal = 16'sd31611;
            8'd212 : out_signal = 16'sd31670;
            8'd213 : out_signal = 16'sd31727;
            8'd214 : out_signal = 16'sd31781;
            8'd215 : out_signal = 16'sd31833;
            8'd216 : out_signal = 16'sd31882;
            8'd217 : out_signal = 16'sd31930;
            8'd218 : out_signal = 16'sd31975;
            8'd219 : out_signal = 16'sd32018;
            8'd220 : out_signal = 16'sd32059;
            8'd221 : out_signal = 16'sd32098;
            8'd222 : out_signal = 16'sd32136;
            8'd223 : out_signal = 16'sd32172;
            8'd224 : out_signal = 16'sd32206;
            8'd225 : out_signal = 16'sd32239;
            8'd226 : out_signal = 16'sd32270;
            8'd227 : out_signal = 16'sd32300;
            8'd228 : out_signal = 16'sd32329;
            8'd229 : out_signal = 16'sd32356;
            8'd230 : out_signal = 16'sd32382;
            8'd231 : out_signal = 16'sd32407;
            8'd232 : out_signal = 16'sd32431;
            8'd233 : out_signal = 16'sd32453;
            8'd234 : out_signal = 16'sd32475;
            8'd235 : out_signal = 16'sd32496;
            8'd236 : out_signal = 16'sd32516;
            8'd237 : out_signal = 16'sd32534;
            8'd238 : out_signal = 16'sd32552;
            8'd239 : out_signal = 16'sd32570;
            8'd240 : out_signal = 16'sd32586;
            8'd241 : out_signal = 16'sd32602;
            8'd242 : out_signal = 16'sd32617;
            8'd243 : out_signal = 16'sd32631;
            8'd244 : out_signal = 16'sd32645;
            8'd245 : out_signal = 16'sd32658;
            8'd246 : out_signal = 16'sd32670;
            8'd247 : out_signal = 16'sd32682;
            8'd248 : out_signal = 16'sd32693;
            8'd249 : out_signal = 16'sd32704;
            8'd250 : out_signal = 16'sd32714;
            8'd251 : out_signal = 16'sd32724;
            8'd252 : out_signal = 16'sd32734;
            8'd253 : out_signal = 16'sd32742;
            8'd254 : out_signal = 16'sd32751;
            8'd255 : out_signal = 16'sd32759;
            default: out_signal = in_signal;
        endcase
    end

endmodule
